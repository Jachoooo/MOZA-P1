* C:\Users\kasia\Desktop\MOZA P1\WSB.asc
RC1 VCC N002 6.8k
RC2 VCC N001 {RC2}
RC3 VCC out 250
RE2 N004 0 {RE2}
Q1 N001 N002 N004 0 2N2222
Q2 out N001 N007 0 2N2222
RE3 N007 0 220
RE1 N005 0 50
CF N006 0 {CF}
RF N006 N005 {RF/2}
RF2 N007 N006 {RF/2}
J1 N002 N003 N005 U309
RS N003 Vin 50
V_AC Vin VDC SINE(0 100m 1k) AC 1
V_DC VDC 0 {VDC}
V_VCC VCC 0 12
.model NPN NPN
.model PNP PNP
.lib C:\Users\kasia\Documents\LTspiceXVII\lib\cmp\standard.bjt
.model NJF NJF
.model PJF PJF
.lib C:\Users\kasia\Documents\LTspiceXVII\lib\cmp\standard.jft
.INCLUDE parametry_inzynierskie.inc
.tran 10m
*.options trtol 5
.backanno
.end
